../kianv_harris_mcycle_edition/gateware/kianv_harris_edition/./riscv_defines.vh